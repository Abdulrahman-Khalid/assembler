LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
library work;

ENTITY EXECUTE_MIR IS 
  PORT(MIR : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
       F1_OUT : OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
       F2_OUT,F3_OUT, F4_OUT,F6_OUT : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
       NEXT_ADDRESS : OUT STD_LOGIC_VECTOR(4 DOWNTO 0));
  END ENTITY EXECUTE_MIR;
  
  
ARCHITECTURE EXECUTE_MIR_ARCH OF EXECUTE_MIR IS
  BEGIN
    F1 : ENTITY WORK.EXECUTE_F1 PORT MAP (MIR(10 DOWNTO 8), F1_OUT);
    F2 : ENTITY WORK.EXECUTE_F2 PORT MAP (MIR(7 DOWNTO 6), F2_OUT);
    F3 : ENTITY WORK.EXECUTE_F3 PORT MAP (MIR(5 DOWNTO 4), F3_OUT);
    F4 : ENTITY WORK.EXECUTE_F4 PORT MAP (MIR(3 DOWNTO 2), F4_OUT); 
    F6 : ENTITY WORK.EXECUTE_F6 PORT MAP (MIR(1 DOWNTO 0), F6_OUT);
    NEXT_ADDRESS <= MIR(15 DOWNTO 11);
   
  END ARCHITECTURE EXECUTE_MIR_ARCH;