LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY EXECUTE_F1 IS
PORT(
  MIR : IN STD_LOGIC_VECTOR( 10 DOWNTO 8);
  EN_TRI_STATE : OUT STD_LOGIC_VECTOR (7 DOWNTO 0)
);

END ENTITY EXECUTE_F1;


ARCHITECTURE EXECUTE_F1_ARCH OF EXECUTE_F1 IS 
BEGIN 
  EN_TRI_STATE <= "00000001" WHEN MIR="000"
             ELSE "00000010" WHEN MIR="001"
             ELSE "00000100" WHEN MIR="010"
             ELSE "00001000" WHEN MIR="011"
             ELSE "00010000" WHEN MIR="100"
             ELSE "00100000" WHEN MIR="101"
             ELSE "01000000" WHEN MIR="110"
             ELSE "10000000" ; 
              
END ARCHITECTURE EXECUTE_F1_ARCH;
