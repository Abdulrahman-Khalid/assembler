LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
library work;

ENTITY ORING IS
  PORT (ENABLE, CLK : IN STD_LOGIC;
        IR : IN STD_LOGIC_VECTOR (15 DOWNTO 0);
        SRC_DEST_SELECTOR : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
        ADRESS : IN STD_LOGIC_VECTOR (15 DOWNTO 11);
        NEXT_ADD : OUT STD_LOGIC_VECTOR (15 DOWNTO 11));

END ENTITY ORING;
  
ARCHITECTURE ORING_ARCH OF ORING IS
  SIGNAL OUT_TWO_OP0, OUT_TWO_OP1, OUT_A2, OUT_B4, OUT_D: STD_LOGIC_VECTOR (15 DOWNTO 11) := "00000";
  SIGNAL EN1, EN2, EN3, EN4, EN5 : STD_LOGIC := '0';
    BEGIN
      
      O1: ENTITY WORK.TWO_OP0_ORING PORT MAP(ENABLE, CLK, IR (15 DOWNTO 12), ADRESS(15 DOWNTO 11), OUT_TWO_OP0(15 DOWNTO 11));  
      O2: ENTITY WORK.TWO_OP1_ORING PORT MAP(ENABLE, CLK, IR (15 DOWNTO 12), ADRESS(15 DOWNTO 11), OUT_TWO_OP1(15 DOWNTO 11));
      O3: ENTITY WORK.A2_ORING PORT MAP (ENABLE, CLK, IR(15 DOWNTO 0),SRC_DEST_SELECTOR, ADRESS(15 DOWNTO 11), OUT_A2(15 DOWNTO 11));
      O4: ENTITY WORK.B4_ORING PORT MAP (ENABLE, CLK, IR(5), IR(11), SRC_DEST_SELECTOR(1 DOWNTO 0), ADRESS(15 DOWNTO 11), OUT_B4(15 DOWNTO 11));
      O5: ENTITY WORK.D_ORING PORT MAP(ENABLE, CLK, IR(14 DOWNTO 6), ADRESS(15 DOWNTO 11) , OUT_D(15 DOWNTO 11));
      
      EN1 <= '1' WHEN ADRESS = "10110" ELSE '0';
      EN2 <= '1' WHEN ADRESS = "10111" ELSE '0';
      EN3 <= '1' WHEN ADRESS = "01010" ELSE '0';
      EN4 <= '1' WHEN ADRESS = "01000" ELSE '0';
      EN5 <= '1' WHEN ADRESS = "01010" ELSE '0';
      
      T1: ENTITY WORK.TRI_STATE PORT MAP (OUT_TWO_OP0(15 DOWNTO 11), EN1, NEXT_ADD(15 DOWNTO 11) );
      T2: ENTITY WORK.TRI_STATE PORT MAP (OUT_TWO_OP1(15 DOWNTO 11), EN2, NEXT_ADD(15 DOWNTO 11) );
      T3: ENTITY WORK.TRI_STATE PORT MAP (OUT_A2(15 DOWNTO 11), EN3, NEXT_ADD(15 DOWNTO 11) );
      T4: ENTITY WORK.TRI_STATE PORT MAP (OUT_B4(15 DOWNTO 11), EN4, NEXT_ADD(15 DOWNTO 11) );
      T5: ENTITY WORK.TRI_STATE PORT MAP (OUT_D(15 DOWNTO 11), EN5, NEXT_ADD(15 DOWNTO 11) ); 
    
      NEXT_ADD <= ADRESS when EN1 = '0' and EN2 = '0' and EN3 = '0' and EN4 = '0' and EN5 = '0';
    
END ARCHITECTURE ORING_ARCH;      
