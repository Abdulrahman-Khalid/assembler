LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
LIBRARY WORK;

ENTITY main IS
	PORT( Clk,Rst : IN std_logic;
	      BUS_DATA	: INOUT   std_logic_vector (15 DOWNTO 0);
		   d : IN std_logic_vector(15 DOWNTO 0);
		   q,qbar : OUT std_logic_vector(15 DOWNTO 0);
		   MIR : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
		   R0 , R1, R2 ,R3, R4, R5, R6, R7 ,DEST, MDR, SRC: INOUT STD_LOGIC_VECTOR (15 DOWNTO 0);
		   MAR : OUT STD_LOGIC_VECTOR (12 DOWNTO 0);
		   RD,WR : OUT STD_LOGIC;
		   IR : IN STD_LOGIC_VECTOR (15 DOWNTO 0));
END main;

ARCHITECTURE main_arch OF main IS
	
	  SIGNAL SEL :STD_LOGIC_VECTOR(1 DOWNTO 0);
	  SIGNAL M_IR :STD_LOGIC_VECTOR(15 DOWNTO 0); 
	  SIGNAL ENAPLE_REGISTER: STD_LOGIC_VECTOR(7 DOWNTO 0);
	  SIGNAL OUT_DEC_SRC,OUT_DEC_DST : STD_LOGIC_VECTOR (7 DOWNTO 0);
	  SIGNAL ADRESS, NEXT_ADDRESS : STD_LOGIC_VECTOR (15 DOWNTO 11);
	  SIGNAL SIG_R0,SIG_R1,SIG_R2,SIG_R3,SIG_R4,SIG_R5,SIG_R6,SIG_R7 : STD_LOGIC_VECTOR (15 DOWNTO 0);
	BEGIN
	   
	    
	   u0: ENTITY WORK.REG GENERIC MAP (16) PORT MAP (BUS_DATA, ENAPLE_REGISTER(0), CLK, RST, R0,qbar);
	   u1: ENTITY WORK.REG GENERIC MAP (16) PORT MAP (BUS_DATA, ENAPLE_REGISTER(1), CLK, RST, R1); 
	   u2: ENTITY WORK.REG GENERIC MAP (16) PORT MAP (BUS_DATA, ENAPLE_REGISTER(2), CLK, RST, R2);
	   u3: ENTITY WORK.REG GENERIC MAP (16) PORT MAP (BUS_DATA, ENAPLE_REGISTER(3), CLK, RST, R3);
	   u4: ENTITY WORK.REG GENERIC MAP (16) PORT MAP (BUS_DATA, ENAPLE_REGISTER(4), CLK, RST, R4);
	   u5: ENTITY WORK.REG GENERIC MAP (16) PORT MAP (BUS_DATA, ENAPLE_REGISTER(5), CLK, RST, R5);
	   u6: ENTITY WORK.REG GENERIC MAP (16) PORT MAP (BUS_DATA, ENAPLE_REGISTER(6), CLK, RST, R6);
	   u7: ENTITY WORK.REG GENERIC MAP (16) PORT MAP (BUS_DATA, ENAPLE_REGISTER(7), CLK, RST, R7);  
 	    
	   
	   OT : ENTITY WORK.OPERATION_TYPE PORT MAP (IR,SEL);
	   FR : ENTITY WORK.FETCH_REGISTERS(IR,R0,R1,R2,R3,R4,R5,R6,R7,SEL,DEST);
	   --FM : ENTITY WORK.FIRST_MIR(IR,SEL,M_IR(15 DOWNTO 11));
	   BD : ENTITY WORK.BIG_DECODER PORT MAP (SEL(1 DOWNTO 0),ADRESS (15 DOWNTO 11), NEXT_ADDRESS(15 DOWNTO 11), IR (15 DOWNTO 0));
	   
	   
	   --DEC_REG_DIR_SRC : DECODER GENERIC MAP (3) PORT MAP (IR(8 DOWNTO 6), OUT_DEC_SRC);
	   --DEC_REG_DIR_DST : DECODER GENERIC MAP (3) PORT MAP (IR(2 DOWNTO 0), OUT_DEC_DST);
	     
    
     --PROCESS
      -- BEGIN
         
       --END PROCESS
	
END main_arch;