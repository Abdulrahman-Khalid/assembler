LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY TWO_OP0_ORING IS
  PORT (IR: IN STD_LOGIC_VECTOR (15 DOWNTO 12);
        ADRESS : IN STD_LOGIC_VECTOR (15 DOWNTO 11);
        NEXT_ADD: OUT STD_LOGIC_VECTOR (15 DOWNTO 11));
    
    
    
END ENTITY TWO_OP0_ORING;
  
ARCHITECTURE TWO_OP0_ORING_ARCH OF TWO_OP0_ORING IS 

BEGIN
  
  NEXT_ADD <= "10111" WHEN ADRESS = "10110" AND IR = "0001" ELSE
              ADRESS;
     
END TWO_OP0_ORING_ARCH;
  
