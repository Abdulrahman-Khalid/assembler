LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
library work;

ENTITY BIG_DECODER IS 
PORT(SRC_DEST_SELECTOR : IN STD_LOGIC_VECTOR (1 DOWNTO 0);
     ADRESS : IN STD_LOGIC_VECTOR ( 15 DOWNTO 11);
     NEXT_ADD : OUT STD_LOGIC_VECTOR ( 15 DOWNTO 11);
     --OUT_NEXT : OUT STD_LOGIC_VECTOR (4 DOWNTO 0);
     IR : IN STD_LOGIC_VECTOR( 15 DOWNTO 0 ));
END ENTITY BIG_DECODER;

ARCHITECTURE BIG_DECODER_ARCH OF BIG_DECODER IS 
SIGNAL NEXT_ADDRESS : STD_LOGIC_VECTOR ( 15 DOWNTO 11); --OUTPUT SIGNAL FROM ORING CIRCUIT AND INPUT TO ROM
SIGNAL MIR : STD_LOGIC_VECTOR (15 DOWNTO 0); --OUTPUT SIGNAL FROM ROM CIRCUIT AND INPUT TO EXECUTE_MIR
SIGNAL F2_OUT1,F3_OUT1, F4_OUT1,F6_OUT1 : STD_LOGIC_VECTOR (3 DOWNTO 0);
SIGNAL F1_OUT1 : STD_LOGIC_VECTOR (7 DOWNTO 0);

BEGIN
  
  O : ENTITY WORK.ORING PORT MAP(IR( 15 DOWNTO 0 ), SRC_DEST_SELECTOR(1 DOWNTO 0), ADRESS(15 DOWNTO 11), NEXT_ADDRESS(15 DOWNTO 11));
  R : ENTITY WORK.ROM PORT MAP(NEXT_ADDRESS(15 DOWNTO 11), MIR( 15 DOWNTO 0));
  E : ENTITY WORK.EXECUTE_MIR PORT MAP(MIR( 15 DOWNTO 0),  F1_OUT1(7 DOWNTO 0), F2_OUT1(3 DOWNTO 0),F3_OUT1(3 DOWNTO 0), F4_OUT1(3 DOWNTO 0),F6_OUT1(3 DOWNTO 0), NEXT_ADD(15 DOWNTO 11));
  
  
END ARCHITECTURE BIG_DECODER_ARCH;  
