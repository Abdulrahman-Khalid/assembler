 LIBRARY IEEE;
USE IEEE.std_logic_1164.all;

ENTITY TWO_OP1_ORING IS
    PORT (IR: IN STD_LOGIC_VECTOR (15 DOWNTO 12);
          ADRESS : IN STD_LOGIC_VECTOR (15 DOWNTO 11);
          NEXT_ADD: OUT STD_LOGIC_VECTOR (15 DOWNTO 11));
         
          
END ENTITY TWO_OP1_ORING;

ARCHITECTURE TWO_OP1_ORING_ARCH OF TWO_OP1_ORING IS
  BEGIN
    
     
  NEXT_ADD <= "00000" WHEN ADRESS = "10111" AND IR = "0010" ELSE
              ADRESS;
    
END ARCHITECTURE TWO_OP1_ORING_ARCH;
  
            
  
